module gen

const (
	main_c = '
int main() {
	v_main_main();
	return 0;
}
'
)