module gen

const (
	std_include = '
#include <default.h>  
'
)