module gen

const (
	std_include = '
#include <stdio.h>  
#include <stdlib.h>
'
)