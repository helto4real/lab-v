module parser

// pub struct Table {
// pub mut:
// 	// types         []TypeSymbol
// 	fns           map[string]Fn
// }

// pub struct Fn {
// pub:
// 	// params         []Param
// 	// return_type    Type
// pub mut:
// 	name      string
// }