module gen

const (
	std_include = '
#include <stdio.h>  
#include <stdlib.h>
#include <stdarg.h> // for va_list
#include <string.h> // memcpy
'
)