module table

pub enum Type {
	string
	unknown
}
