module gen

const (
	std_include = '
#include <stdio.h>  // TODO remove all these includes, define all function signatures and types manually
#include <stdlib.h>
'
)